//                              -*- Mode: Verilog -*-
// Filename        : ipcore.sv
// Description     : Example ipcore
// Author          : Adrian Fiergolski
// Created On      : Thu Sep 18 11:00:12 2014
// Last Modified By: Adrian Fiergolski
// Last Modified On: Thu Sep 18 11:00:12 2014
// Update Count    : 0
// Status          : Unknown, Use with caution!

`include "ipcoreInclude.sv"

module ipcore;
   ipcoreInclude incl();
endmodule // ipcore
