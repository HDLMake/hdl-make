//                              -*- Mode: Verilog -*-
// Filename        : ipcoreInclude.sv
// Description     : Example ipcoreinclude
// Author          : Adrian Fiergolski
// Created On      : Thu Sep 18 11:01:31 2014
// Last Modified By: Adrian Fiergolski
// Last Modified On: Thu Sep 18 11:01:31 2014
// Update Count    : 0
// Status          : Unknown, Use with caution!

module ipcoreInclude;
endmodule // ipcoreinclude
