-- This file has been generated with Libre-FDATool
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.all;

ENTITY tb_myfilter IS
END tb_myfilter;

ARCHITECTURE behavior OF tb_myfilter IS
    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT myfilter
    PORT(
        clk: IN std_logic;
        rst: IN std_logic;
        sig_in: IN signed(15 downto 0);
        sig_out: OUT signed(15 downto 0)
    );
    END COMPONENT;

    -- Signal Declaration
    signal clk : std_logic := '0';
    signal rst : std_logic := '1';
    signal sig_in : signed(15 downto 0);
    signal sig_out : signed(15 downto 0);

BEGIN
    -- Instantiate the Unit Under Test (UUT)
    uut: myfilter PORT MAP (
        clk => clk,
        rst => rst,
        sig_in => sig_in,
        sig_out => sig_out
    );

    clk_process : process
    begin
        clk <= '1';
        wait for 25 ns;
        clk <= '0';
        wait for 25 ns;
    end process;
    stimulus_process : process
    begin
        sig_in <=  (others => '0');
        rst <= '1'; wait for 100 ns;
        rst <= '0'; wait for 125 ns;
        wait for 50 ns; sig_in <= "0000000000000000"; -- -0.000000
        wait for 50 ns; sig_in <= "0000000000000101"; -- 0.000157
        wait for 50 ns; sig_in <= "0000000000010101"; -- 0.000630
        wait for 50 ns; sig_in <= "0000000000101110"; -- 0.001417
        wait for 50 ns; sig_in <= "0000000001010011"; -- 0.002518
        wait for 50 ns; sig_in <= "0000000010000001"; -- 0.003935
        wait for 50 ns; sig_in <= "0000000010111010"; -- 0.005666
        wait for 50 ns; sig_in <= "0000000011111101"; -- 0.007712
        wait for 50 ns; sig_in <= "0000000101001010"; -- 0.010073
        wait for 50 ns; sig_in <= "0000000110100010"; -- 0.012748
        wait for 50 ns; sig_in <= "0000001000000100"; -- 0.015737
        wait for 50 ns; sig_in <= "0000001001110000"; -- 0.019040
        wait for 50 ns; sig_in <= "0000001011100110"; -- 0.022657
        wait for 50 ns; sig_in <= "0000001101100111"; -- 0.026587
        wait for 50 ns; sig_in <= "0000001111110010"; -- 0.030830
        wait for 50 ns; sig_in <= "0000010010000111"; -- 0.035384
        wait for 50 ns; sig_in <= "0000010100100111"; -- 0.040249
        wait for 50 ns; sig_in <= "0000010111010000"; -- 0.045424
        wait for 50 ns; sig_in <= "0000011010000100"; -- 0.050907
        wait for 50 ns; sig_in <= "0000011101000010"; -- 0.056697
        wait for 50 ns; sig_in <= "0000100000001010"; -- 0.062791
        wait for 50 ns; sig_in <= "0000100011011011"; -- 0.069188
        wait for 50 ns; sig_in <= "0000100110110111"; -- 0.075884
        wait for 50 ns; sig_in <= "0000101010011100"; -- 0.082877
        wait for 50 ns; sig_in <= "0000101110001010"; -- 0.090163
        wait for 50 ns; sig_in <= "0000110010000011"; -- 0.097738
        wait for 50 ns; sig_in <= "0000110110000100"; -- 0.105597
        wait for 50 ns; sig_in <= "0000111010001111"; -- 0.113736
        wait for 50 ns; sig_in <= "0000111110100011"; -- 0.122148
        wait for 50 ns; sig_in <= "0001000010111111"; -- 0.130828
        wait for 50 ns; sig_in <= "0001000111100100"; -- 0.139767
        wait for 50 ns; sig_in <= "0001001100010001"; -- 0.148959
        wait for 50 ns; sig_in <= "0001010001000110"; -- 0.158395
        wait for 50 ns; sig_in <= "0001010110000011"; -- 0.168065
        wait for 50 ns; sig_in <= "0001011011000111"; -- 0.177959
        wait for 50 ns; sig_in <= "0001100000010011"; -- 0.188065
        wait for 50 ns; sig_in <= "0001100101100100"; -- 0.198372
        wait for 50 ns; sig_in <= "0001101010111100"; -- 0.208865
        wait for 50 ns; sig_in <= "0001110000011010"; -- 0.219531
        wait for 50 ns; sig_in <= "0001110101111100"; -- 0.230354
        wait for 50 ns; sig_in <= "0001111011100100"; -- 0.241318
        wait for 50 ns; sig_in <= "0010000001001111"; -- 0.252404
        wait for 50 ns; sig_in <= "0010000110111101"; -- 0.263594
        wait for 50 ns; sig_in <= "0010001100101111"; -- 0.274866
        wait for 50 ns; sig_in <= "0010010010100010"; -- 0.286200
        wait for 50 ns; sig_in <= "0010011000010111"; -- 0.297573
        wait for 50 ns; sig_in <= "0010011110001100"; -- 0.308959
        wait for 50 ns; sig_in <= "0010100100000001"; -- 0.320334
        wait for 50 ns; sig_in <= "0010101001110100"; -- 0.331670
        wait for 50 ns; sig_in <= "0010101111100101"; -- 0.342938
        wait for 50 ns; sig_in <= "0010110101010011"; -- 0.354109
        wait for 50 ns; sig_in <= "0010111010111101"; -- 0.365151
        wait for 50 ns; sig_in <= "0011000000100010"; -- 0.376032
        wait for 50 ns; sig_in <= "0011000110000000"; -- 0.386717
        wait for 50 ns; sig_in <= "0011001011010110"; -- 0.397171
        wait for 50 ns; sig_in <= "0011010000100100"; -- 0.407357
        wait for 50 ns; sig_in <= "0011010101101000"; -- 0.417237
        wait for 50 ns; sig_in <= "0011011010100000"; -- 0.426771
        wait for 50 ns; sig_in <= "0011011111001100"; -- 0.435921
        wait for 50 ns; sig_in <= "0011100011101010"; -- 0.444642
        wait for 50 ns; sig_in <= "0011100111111000"; -- 0.452895
        wait for 50 ns; sig_in <= "0011101011110110"; -- 0.460634
        wait for 50 ns; sig_in <= "0011101111100001"; -- 0.467816
        wait for 50 ns; sig_in <= "0011110010111001"; -- 0.474397
        wait for 50 ns; sig_in <= "0011110101111011"; -- 0.480331
        wait for 50 ns; sig_in <= "0011111000100111"; -- 0.485572
        wait for 50 ns; sig_in <= "0011111010111011"; -- 0.490075
        wait for 50 ns; sig_in <= "0011111100110101"; -- 0.493795
        wait for 50 ns; sig_in <= "0011111110010011"; -- 0.496685
        wait for 50 ns; sig_in <= "0011111111010101"; -- 0.498701
        wait for 50 ns; sig_in <= "0011111111111001"; -- 0.499799
        wait for 50 ns; sig_in <= "0011111111111110"; -- 0.499936
        wait for 50 ns; sig_in <= "0011111111100001"; -- 0.499068
        wait for 50 ns; sig_in <= "0011111110100011"; -- 0.497156
        wait for 50 ns; sig_in <= "0011111101000001"; -- 0.494160
        wait for 50 ns; sig_in <= "0011111010111010"; -- 0.490044
        wait for 50 ns; sig_in <= "0011111000001101"; -- 0.484773
        wait for 50 ns; sig_in <= "0011110100111001"; -- 0.478316
        wait for 50 ns; sig_in <= "0011110000111110"; -- 0.470643
        wait for 50 ns; sig_in <= "0011101100011010"; -- 0.461729
        wait for 50 ns; sig_in <= "0011100111001100"; -- 0.451552
        wait for 50 ns; sig_in <= "0011100001010101"; -- 0.440096
        wait for 50 ns; sig_in <= "0011011010110011"; -- 0.427345
        wait for 50 ns; sig_in <= "0011010011100111"; -- 0.413293
        wait for 50 ns; sig_in <= "0011001011110000"; -- 0.397936
        wait for 50 ns; sig_in <= "0011000011001110"; -- 0.381275
        wait for 50 ns; sig_in <= "0010111010000001"; -- 0.363319
        wait for 50 ns; sig_in <= "0010110000001011"; -- 0.344083
        wait for 50 ns; sig_in <= "0010100101101011"; -- 0.323587
        wait for 50 ns; sig_in <= "0010011010100011"; -- 0.301857
        wait for 50 ns; sig_in <= "0010001110110100"; -- 0.278930
        wait for 50 ns; sig_in <= "0010000010011111"; -- 0.254847
        wait for 50 ns; sig_in <= "0001110101100101"; -- 0.229657
        wait for 50 ns; sig_in <= "0001101000001010"; -- 0.203417
        wait for 50 ns; sig_in <= "0001011010001110"; -- 0.176194
        wait for 50 ns; sig_in <= "0001001011110100"; -- 0.148059
        wait for 50 ns; sig_in <= "0000111100111111"; -- 0.119095
        wait for 50 ns; sig_in <= "0000101101110001"; -- 0.089391
        wait for 50 ns; sig_in <= "0000011110001111"; -- 0.059044
        wait for 50 ns; sig_in <= "0000001110011011"; -- 0.028160
        wait for 50 ns; sig_in <= "1111111110011001"; -- -0.003146
        wait for 50 ns; sig_in <= "1111101110001101"; -- -0.034755
        wait for 50 ns; sig_in <= "1111011101111100"; -- -0.066536
        wait for 50 ns; sig_in <= "1111001101101001"; -- -0.098354
        wait for 50 ns; sig_in <= "1110111101011010"; -- -0.130067
        wait for 50 ns; sig_in <= "1110101101010011"; -- -0.161525
        wait for 50 ns; sig_in <= "1110011101011010"; -- -0.192575
        wait for 50 ns; sig_in <= "1110001101110011"; -- -0.223058
        wait for 50 ns; sig_in <= "1101111110100100"; -- -0.252810
        wait for 50 ns; sig_in <= "1101101111110010"; -- -0.281665
        wait for 50 ns; sig_in <= "1101100001100100"; -- -0.309453
        wait for 50 ns; sig_in <= "1101010011111110"; -- -0.336004
        wait for 50 ns; sig_in <= "1101000111000110"; -- -0.361147
        wait for 50 ns; sig_in <= "1100111011000010"; -- -0.384713
        wait for 50 ns; sig_in <= "1100101111110111"; -- -0.406533
        wait for 50 ns; sig_in <= "1100100101101010"; -- -0.426442
        wait for 50 ns; sig_in <= "1100011100100010"; -- -0.444281
        wait for 50 ns; sig_in <= "1100010100100010"; -- -0.459895
        wait for 50 ns; sig_in <= "1100001101110000"; -- -0.473139
        wait for 50 ns; sig_in <= "1100001000010000"; -- -0.483873
        wait for 50 ns; sig_in <= "1100000100000111"; -- -0.491972
        wait for 50 ns; sig_in <= "1100000001011000"; -- -0.497321
        wait for 50 ns; sig_in <= "1100000000000110"; -- -0.499817
        wait for 50 ns; sig_in <= "1100000000010101"; -- -0.499374
        wait for 50 ns; sig_in <= "1100000010000110"; -- -0.495922
        wait for 50 ns; sig_in <= "1100000101011011"; -- -0.489410
        wait for 50 ns; sig_in <= "1100001010010110"; -- -0.479804
        wait for 50 ns; sig_in <= "1100010000110110"; -- -0.467091
        wait for 50 ns; sig_in <= "1100011000111100"; -- -0.451282
        wait for 50 ns; sig_in <= "1100100010100111"; -- -0.432409
        wait for 50 ns; sig_in <= "1100101101110100"; -- -0.410528
        wait for 50 ns; sig_in <= "1100111010100001"; -- -0.385719
        wait for 50 ns; sig_in <= "1101001000101010"; -- -0.358089
        wait for 50 ns; sig_in <= "1101011000001100"; -- -0.327768
        wait for 50 ns; sig_in <= "1101101001000000"; -- -0.294913
        wait for 50 ns; sig_in <= "1101111011000010"; -- -0.259707
        wait for 50 ns; sig_in <= "1110001110001010"; -- -0.222358
        wait for 50 ns; sig_in <= "1110100010010000"; -- -0.183099
        wait for 50 ns; sig_in <= "1110110111001101"; -- -0.142187
        wait for 50 ns; sig_in <= "1111001100110110"; -- -0.099901
        wait for 50 ns; sig_in <= "1111100011000011"; -- -0.056544
        wait for 50 ns; sig_in <= "1111111001101000"; -- -0.012436
        wait for 50 ns; sig_in <= "0000010000011011"; -- 0.032083
        wait for 50 ns; sig_in <= "0000100111010000"; -- 0.076659
        wait for 50 ns; sig_in <= "0000111101111010"; -- 0.120924
        wait for 50 ns; sig_in <= "0001010100001110"; -- 0.164500
        wait for 50 ns; sig_in <= "0001101001111111"; -- 0.207001
        wait for 50 ns; sig_in <= "0001111111000000"; -- 0.248041
        wait for 50 ns; sig_in <= "0010010011000100"; -- 0.287229
        wait for 50 ns; sig_in <= "0010100101111111"; -- 0.324182
        wait for 50 ns; sig_in <= "0010110111100100"; -- 0.358524
        wait for 50 ns; sig_in <= "0011000111101000"; -- 0.389888
        wait for 50 ns; sig_in <= "0011010101111111"; -- 0.417928
        wait for 50 ns; sig_in <= "0011100010011110"; -- 0.442315
        wait for 50 ns; sig_in <= "0011101100111011"; -- 0.462747
        wait for 50 ns; sig_in <= "0011110101001110"; -- 0.478952
        wait for 50 ns; sig_in <= "0011111011001111"; -- 0.490689
        wait for 50 ns; sig_in <= "0011111110110110"; -- 0.497757
        wait for 50 ns; sig_in <= "0100000000000000"; -- 0.499995
        wait for 50 ns; sig_in <= "0011111110100111"; -- 0.497289
        wait for 50 ns; sig_in <= "0011111010101010"; -- 0.489571
        wait for 50 ns; sig_in <= "0011110100001001"; -- 0.476826
        wait for 50 ns; sig_in <= "0011101011000100"; -- 0.459091
        wait for 50 ns; sig_in <= "0011011111011110"; -- 0.436461
        wait for 50 ns; sig_in <= "0011010001011101"; -- 0.409086
        wait for 50 ns; sig_in <= "0011000001000111"; -- 0.377174
        wait for 50 ns; sig_in <= "0010101110100110"; -- 0.340990
        wait for 50 ns; sig_in <= "0010011010000010"; -- 0.300855
        wait for 50 ns; sig_in <= "0010000011101010"; -- 0.257148
        wait for 50 ns; sig_in <= "0001101011101011"; -- 0.210298
        wait for 50 ns; sig_in <= "0001010010010101"; -- 0.160786
        wait for 50 ns; sig_in <= "0000110111111000"; -- 0.109138
        wait for 50 ns; sig_in <= "0000011100101000"; -- 0.055920
        wait for 50 ns; sig_in <= "0000000000111001"; -- 0.001736
        wait for 50 ns; sig_in <= "1111100100111110"; -- -0.052781
        wait for 50 ns; sig_in <= "1111001001001111"; -- -0.106977
        wait for 50 ns; sig_in <= "1110101101111111"; -- -0.160181
        wait for 50 ns; sig_in <= "1110010011100110"; -- -0.211717
        wait for 50 ns; sig_in <= "1101111010011011"; -- -0.260909
        wait for 50 ns; sig_in <= "1101100010110001"; -- -0.307096
        wait for 50 ns; sig_in <= "1101001100111111"; -- -0.349633
        wait for 50 ns; sig_in <= "1100111001011001"; -- -0.387909
        wait for 50 ns; sig_in <= "1100101000010001"; -- -0.421350
        wait for 50 ns; sig_in <= "1100011001111001"; -- -0.449433
        wait for 50 ns; sig_in <= "1100001110100000"; -- -0.471694
        wait for 50 ns; sig_in <= "1100000110010010"; -- -0.487736
        wait for 50 ns; sig_in <= "1100000001011010"; -- -0.497238
        wait for 50 ns; sig_in <= "1100000000000001"; -- -0.499962
        wait for 50 ns; sig_in <= "1100000010001011"; -- -0.495761
        wait for 50 ns; sig_in <= "1100000111111001"; -- -0.484581
        wait for 50 ns; sig_in <= "1100010001001011"; -- -0.466472
        wait for 50 ns; sig_in <= "1100011101111010"; -- -0.441583
        wait for 50 ns; sig_in <= "1100101110000000"; -- -0.410170
        wait for 50 ns; sig_in <= "1101000001001111"; -- -0.372593
        wait for 50 ns; sig_in <= "1101010111011001"; -- -0.329312
        wait for 50 ns; sig_in <= "1101110000001100"; -- -0.280890
        wait for 50 ns; sig_in <= "1110001011010001"; -- -0.227982
        wait for 50 ns; sig_in <= "1110101000010010"; -- -0.171328
        wait for 50 ns; sig_in <= "1111000110110010"; -- -0.111749
        wait for 50 ns; sig_in <= "1111100110010101"; -- -0.050131
        wait for 50 ns; sig_in <= "0000000110011100"; -- 0.012584
        wait for 50 ns; sig_in <= "0000100110100111"; -- 0.075411
        wait for 50 ns; sig_in <= "0001000110010100"; -- 0.137342
        wait for 50 ns; sig_in <= "0001100101000011"; -- 0.197354
        wait for 50 ns; sig_in <= "0010000010010001"; -- 0.254434
        wait for 50 ns; sig_in <= "0010011101011111"; -- 0.307591
        wait for 50 ns; sig_in <= "0010110110001101"; -- 0.355878
        wait for 50 ns; sig_in <= "0011001011111111"; -- 0.398407
        wait for 50 ns; sig_in <= "0011011110011001"; -- 0.434367
        wait for 50 ns; sig_in <= "0011101101000101"; -- 0.463044
        wait for 50 ns; sig_in <= "0011110111101110"; -- 0.483833
        wait for 50 ns; sig_in <= "0011111110000101"; -- 0.496255
        wait for 50 ns; sig_in <= "0011111111111111"; -- 0.499971
        wait for 50 ns; sig_in <= "0011111101010101"; -- 0.494791
        wait for 50 ns; sig_in <= "0011110110000111"; -- 0.480681
        wait for 50 ns; sig_in <= "0011101010011000"; -- 0.457773
        wait for 50 ns; sig_in <= "0011011010010011"; -- 0.426365
        wait for 50 ns; sig_in <= "0011000110000111"; -- 0.386921
        wait for 50 ns; sig_in <= "0010101110000111"; -- 0.340070
        wait for 50 ns; sig_in <= "0010010010101111"; -- 0.286594
        wait for 50 ns; sig_in <= "0001110100011100"; -- 0.227423
        wait for 50 ns; sig_in <= "0001010011110001"; -- 0.163618
        wait for 50 ns; sig_in <= "0000110001010101"; -- 0.096356
        wait for 50 ns; sig_in <= "0000001101110010"; -- 0.026909
        wait for 50 ns; sig_in <= "1111101001110011"; -- -0.043378
        wait for 50 ns; sig_in <= "1111000110000101"; -- -0.113115
        wait for 50 ns; sig_in <= "1110100011011001"; -- -0.180890
        wait for 50 ns; sig_in <= "1110000010011010"; -- -0.245299
        wait for 50 ns; sig_in <= "1101100011110111"; -- -0.304977
        wait for 50 ns; sig_in <= "1101001000011000"; -- -0.358630
        wait for 50 ns; sig_in <= "1100110000100111"; -- -0.405058
        wait for 50 ns; sig_in <= "1100011101000110"; -- -0.443190
        wait for 50 ns; sig_in <= "1100001110010010"; -- -0.472109
        wait for 50 ns; sig_in <= "1100000100100100"; -- -0.491077
        wait for 50 ns; sig_in <= "1100000000001111"; -- -0.499555
        wait for 50 ns; sig_in <= "1100000001011011"; -- -0.497223
        wait for 50 ns; sig_in <= "1100001000001100"; -- -0.483995
        wait for 50 ns; sig_in <= "1100010100011110"; -- -0.460023
        wait for 50 ns; sig_in <= "1100100110000010"; -- -0.425707
        wait for 50 ns; sig_in <= "1100111100100101"; -- -0.381687
        wait for 50 ns; sig_in <= "1101010111101001"; -- -0.328841
        wait for 50 ns; sig_in <= "1101110110101001"; -- -0.268267
        wait for 50 ns; sig_in <= "1110011000111101"; -- -0.201266
        wait for 50 ns; sig_in <= "1110111101110011"; -- -0.129317
        wait for 50 ns; sig_in <= "1111100100010101"; -- -0.054047
        wait for 50 ns; sig_in <= "0000001011101011"; -- 0.022805
        wait for 50 ns; sig_in <= "0000110010111010"; -- 0.099426
        wait for 50 ns; sig_in <= "0001011001000101"; -- 0.173972
        wait for 50 ns; sig_in <= "0001111101001111"; -- 0.244611
        wait for 50 ns; sig_in <= "0010011110100000"; -- 0.309570
        wait for 50 ns; sig_in <= "0010111100000000"; -- 0.367181
        wait for 50 ns; sig_in <= "0011010100111101"; -- 0.415926
        wait for 50 ns; sig_in <= "0011101000101100"; -- 0.454478
        wait for 50 ns; sig_in <= "0011110110101010"; -- 0.481745
        wait for 50 ns; sig_in <= "0011111110011010"; -- 0.496898
        wait for 50 ns; sig_in <= "0011111111101101"; -- 0.499405
        wait for 50 ns; sig_in <= "0011111010011001"; -- 0.489054
        wait for 50 ns; sig_in <= "0011101110100101"; -- 0.465962
        wait for 50 ns; sig_in <= "0011011100011101"; -- 0.430585
        wait for 50 ns; sig_in <= "0011000100011110"; -- 0.383714
        wait for 50 ns; sig_in <= "0010100111001010"; -- 0.326464
        wait for 50 ns; sig_in <= "0010000101010000"; -- 0.260251
        wait for 50 ns; sig_in <= "0001011111101000"; -- 0.186762
        wait for 50 ns; sig_in <= "0000110111010000"; -- 0.107915
        wait for 50 ns; sig_in <= "0000001101001110"; -- 0.025812
        wait for 50 ns; sig_in <= "1111100010101010"; -- -0.057312
        wait for 50 ns; sig_in <= "1110111000110000"; -- -0.139152
        wait for 50 ns; sig_in <= "1110010000101100"; -- -0.217398
        wait for 50 ns; sig_in <= "1101101011101000"; -- -0.289794
        wait for 50 ns; sig_in <= "1101001010101001"; -- -0.354212
        wait for 50 ns; sig_in <= "1100101110101111"; -- -0.408715
        wait for 50 ns; sig_in <= "1100011000110001"; -- -0.451615
        wait for 50 ns; sig_in <= "1100001001011101"; -- -0.481533
        wait for 50 ns; sig_in <= "1100000001010100"; -- -0.497448
        wait for 50 ns; sig_in <= "1100000000101001"; -- -0.498736
        wait for 50 ns; sig_in <= "1100000111100101"; -- -0.485197
        wait for 50 ns; sig_in <= "1100010101111111"; -- -0.457076
        wait for 50 ns; sig_in <= "1100101011011111"; -- -0.415063
        wait for 50 ns; sig_in <= "1101000111100010"; -- -0.360285
        wait for 50 ns; sig_in <= "1101101001010101"; -- -0.294284
        wait for 50 ns; sig_in <= "1110001111111001"; -- -0.218977
        wait for 50 ns; sig_in <= "1110111010000100"; -- -0.136603
        wait for 50 ns; sig_in <= "1111100110100101"; -- -0.049667
        wait for 50 ns; sig_in <= "0000010100000010"; -- 0.039139
        wait for 50 ns; sig_in <= "0001000001000010"; -- 0.127014
        wait for 50 ns; sig_in <= "0001101100000111"; -- 0.211139
        wait for 50 ns; sig_in <= "0010010011110110"; -- 0.288766
        wait for 50 ns; sig_in <= "0010110110111100"; -- 0.357308
        wait for 50 ns; sig_in <= "0011010100001100"; -- 0.414433
        wait for 50 ns; sig_in <= "0011101010100100"; -- 0.458144
        wait for 50 ns; sig_in <= "0011111001010001"; -- 0.486853
        wait for 50 ns; sig_in <= "0011111111101110"; -- 0.499449
        wait for 50 ns; sig_in <= "0011111101100111"; -- 0.495343
        wait for 50 ns; sig_in <= "0011110010111100"; -- 0.474501
        wait for 50 ns; sig_in <= "0011011111111111"; -- 0.437461
        wait for 50 ns; sig_in <= "0011000101010010"; -- 0.385326
        wait for 50 ns; sig_in <= "0010100011101101"; -- 0.319740
        wait for 50 ns; sig_in <= "0001111100010110"; -- 0.242845
        wait for 50 ns; sig_in <= "0001010000100000"; -- 0.157214
        wait for 50 ns; sig_in <= "0000100001101011"; -- 0.065771
        wait for 50 ns; sig_in <= "1111110001100001"; -- -0.028302
        wait for 50 ns; sig_in <= "1111000001101101"; -- -0.121677
        wait for 50 ns; sig_in <= "1110010011111110"; -- -0.210995
        wait for 50 ns; sig_in <= "1101101001111111"; -- -0.292989
        wait for 50 ns; sig_in <= "1101000101010101"; -- -0.364604
        wait for 50 ns; sig_in <= "1100100111010111"; -- -0.423115
        wait for 50 ns; sig_in <= "1100010001010010"; -- -0.466237
        wait for 50 ns; sig_in <= "1100000011111111"; -- -0.492221
        wait for 50 ns; sig_in <= "1100000000000010"; -- -0.499928
        wait for 50 ns; sig_in <= "1100000101101100"; -- -0.488891
        wait for 50 ns; sig_in <= "1100010100110100"; -- -0.459345
        wait for 50 ns; sig_in <= "1100101100111100"; -- -0.412235
        wait for 50 ns; sig_in <= "1101001101001110"; -- -0.349197
        wait for 50 ns; sig_in <= "1101110100011110"; -- -0.272508
        wait for 50 ns; sig_in <= "1110100001010001"; -- -0.185013
        wait for 50 ns; sig_in <= "1111010001111010"; -- -0.090024
        wait for 50 ns; sig_in <= "0000000100100000"; -- 0.008798
        wait for 50 ns; sig_in <= "0000110111000101"; -- 0.107581
        wait for 50 ns; sig_in <= "0001100111101000"; -- 0.202395
        wait for 50 ns; sig_in <= "0010010100001011"; -- 0.289405
        wait for 50 ns; sig_in <= "0010111010111001"; -- 0.365033
        wait for 50 ns; sig_in <= "0011011010001011"; -- 0.426106
        wait for 50 ns; sig_in <= "0011110000101001"; -- 0.469996
        wait for 50 ns; sig_in <= "0011111101010100"; -- 0.494742
        wait for 50 ns; sig_in <= "0011111111100100"; -- 0.499144
        wait for 50 ns; sig_in <= "0011110111001101"; -- 0.482831
        wait for 50 ns; sig_in <= "0011100100100000"; -- 0.446294
        wait for 50 ns; sig_in <= "0011001000001000"; -- 0.390884
        wait for 50 ns; sig_in <= "0010100011001110"; -- 0.318774
        wait for 50 ns; sig_in <= "0001110111001111"; -- 0.232880
        wait for 50 ns; sig_in <= "0001000110000001"; -- 0.136759
        wait for 50 ns; sig_in <= "0000010001101001"; -- 0.034459
        wait for 50 ns; sig_in <= "1111011100010110"; -- -0.069639
        wait for 50 ns; sig_in <= "1110101000011100"; -- -0.171010
        wait for 50 ns; sig_in <= "1101111000001111"; -- -0.265182
        wait for 50 ns; sig_in <= "1101001101110111"; -- -0.347932
        wait for 50 ns; sig_in <= "1100101011010001"; -- -0.415484
        wait for 50 ns; sig_in <= "1100010010000101"; -- -0.464684
        wait for 50 ns; sig_in <= "1100000011100000"; -- -0.493159
        wait for 50 ns; sig_in <= "1100000000010010"; -- -0.499436
        wait for 50 ns; sig_in <= "1100001000101100"; -- -0.483035
        wait for 50 ns; sig_in <= "1100011100011010"; -- -0.444507
        wait for 50 ns; sig_in <= "1100111010101010"; -- -0.385429
        wait for 50 ns; sig_in <= "1101100010001000"; -- -0.308355
        wait for 50 ns; sig_in <= "1110010001000011"; -- -0.216716
        wait for 50 ns; sig_in <= "1111000101010010"; -- -0.114674
        wait for 50 ns; sig_in <= "1111111100011100"; -- -0.006944
        wait for 50 ns; sig_in <= "0000110011111011"; -- 0.101421
        wait for 50 ns; sig_in <= "0001101001000110"; -- 0.205266
        wait for 50 ns; sig_in <= "0010011001011001"; -- 0.299578
        wait for 50 ns; sig_in <= "0011000010011011"; -- 0.379730
        wait for 50 ns; sig_in <= "0011100010001010"; -- 0.441719
        wait for 50 ns; sig_in <= "0011110110111110"; -- 0.482369
        wait for 50 ns; sig_in <= "0011111111110000"; -- 0.499507
        wait for 50 ns; sig_in <= "0011111011111101"; -- 0.492088
        wait for 50 ns; sig_in <= "0011101011101010"; -- 0.460274
        wait for 50 ns; sig_in <= "0011001111100110"; -- 0.405443
        wait for 50 ns; sig_in <= "0010101001000010"; -- 0.330151
        wait for 50 ns; sig_in <= "0001111001110111"; -- 0.238021
        wait for 50 ns; sig_in <= "0001000100011001"; -- 0.133580
        wait for 50 ns; sig_in <= "0000001011010010"; -- 0.022049
        wait for 50 ns; sig_in <= "1111010001011101"; -- -0.090917
        wait for 50 ns; sig_in <= "1110011001110111"; -- -0.199508
        wait for 50 ns; sig_in <= "1101100111011001"; -- -0.298062
        wait for 50 ns; sig_in <= "1100111100110000"; -- -0.381362
        wait for 50 ns; sig_in <= "1100011100001101"; -- -0.444921
        wait for 50 ns; sig_in <= "1100000111100100"; -- -0.485227
        wait for 50 ns; sig_in <= "1100000000000001"; -- -0.499958
        wait for 50 ns; sig_in <= "1100000110000101"; -- -0.488120
        wait for 50 ns; sig_in <= "1100011001100010"; -- -0.450132
        wait for 50 ns; sig_in <= "1100111001011100"; -- -0.387826
        wait for 50 ns; sig_in <= "1101100100001010"; -- -0.304377
        wait for 50 ns; sig_in <= "1110010111011110"; -- -0.204155
        wait for 50 ns; sig_in <= "1111010000101001"; -- -0.092506
        wait for 50 ns; sig_in <= "0000001100100100"; -- 0.024522
        wait for 50 ns; sig_in <= "0001000111111100"; -- 0.140502
        wait for 50 ns; sig_in <= "0001111111011111"; -- 0.248980
        wait for 50 ns; sig_in <= "0010110000000011"; -- 0.343837
        wait for 50 ns; sig_in <= "0011010110110111"; -- 0.419637
        wait for 50 ns; sig_in <= "0011110001101001"; -- 0.471949
        wait for 50 ns; sig_in <= "0011111110110010"; -- 0.497619
        wait for 50 ns; sig_in <= "0011111101011011"; -- 0.494973
        wait for 50 ns; sig_in <= "0011101101100010"; -- 0.463940
        wait for 50 ns; sig_in <= "0011001111111011"; -- 0.406089
        wait for 50 ns; sig_in <= "0010100110001011"; -- 0.324562
        wait for 50 ns; sig_in <= "0001110010101010"; -- 0.223925
        wait for 50 ns; sig_in <= "0000111000010010"; -- 0.109924
        wait for 50 ns; sig_in <= "1111111010011101"; -- -0.010836
        wait for 50 ns; sig_in <= "1110111100110011"; -- -0.131261
        wait for 50 ns; sig_in <= "1110000010111110"; -- -0.244187
        wait for 50 ns; sig_in <= "1101010000011111"; -- -0.342806
        wait for 50 ns; sig_in <= "1100101000011010"; -- -0.421085
        wait for 50 ns; sig_in <= "1100001101001111"; -- -0.474140
        wait for 50 ns; sig_in <= "1100000000101111"; -- -0.498560
        wait for 50 ns; sig_in <= "1100000011110001"; -- -0.492637
        wait for 50 ns; sig_in <= "1100010110010001"; -- -0.456505
        wait for 50 ns; sig_in <= "1100110111001110"; -- -0.392162
        wait for 50 ns; sig_in <= "1101100100101011"; -- -0.303380
        wait for 50 ns; sig_in <= "1110011011111010"; -- -0.195501
        wait for 50 ns; sig_in <= "1111011001100010"; -- -0.075131
        wait for 50 ns; sig_in <= "0000011001101111"; -- 0.050256
        wait for 50 ns; sig_in <= "0001011000011110"; -- 0.172776
        wait for 50 ns; sig_in <= "0010010001101111"; -- 0.284629
        wait for 50 ns; sig_in <= "0011000001110110"; -- 0.378597
        wait for 50 ns; sig_in <= "0011100101101001"; -- 0.448524
        wait for 50 ns; sig_in <= "0011111010101111"; -- 0.489724
        wait for 50 ns; sig_in <= "0011111111101010"; -- 0.499319
        wait for 50 ns; sig_in <= "0011110011111100"; -- 0.476452
        wait for 50 ns; sig_in <= "0011011000010001"; -- 0.422380
        wait for 50 ns; sig_in <= "0010101110010011"; -- 0.340430
        wait for 50 ns; sig_in <= "0001111000101111"; -- 0.235808
        wait for 50 ns; sig_in <= "0000111011000010"; -- 0.115294
        wait for 50 ns; sig_in <= "1111111001010000"; -- -0.013193
        wait for 50 ns; sig_in <= "1110110111110000"; -- -0.141101
        wait for 50 ns; sig_in <= "1101111010111110"; -- -0.259816
        wait for 50 ns; sig_in <= "1101000111000011"; -- -0.361239
        wait for 50 ns; sig_in <= "1100011111100100"; -- -0.438352
        wait for 50 ns; sig_in <= "1100000111010100"; -- -0.485715
        wait for 50 ns; sig_in <= "1100000000000100"; -- -0.499865
        wait for 50 ns; sig_in <= "1100001010011101"; -- -0.479589
        wait for 50 ns; sig_in <= "1100100101110111"; -- -0.426047
        wait for 50 ns; sig_in <= "1101010000100001"; -- -0.342730
        wait for 50 ns; sig_in <= "1110000111100011"; -- -0.235255
        wait for 50 ns; sig_in <= "1111000111001011"; -- -0.111003
        wait for 50 ns; sig_in <= "0000001010111100"; -- 0.021371
        wait for 50 ns; sig_in <= "0001001110000110"; -- 0.152534
        wait for 50 ns; sig_in <= "0010001011110110"; -- 0.273131
        wait for 50 ns; sig_in <= "0010111111101110"; -- 0.374453
        wait for 50 ns; sig_in <= "0011100101111011"; -- 0.449077
        wait for 50 ns; sig_in <= "0011111011100111"; -- 0.491425
        wait for 50 ns; sig_in <= "0011111111000101"; -- 0.498198
        wait for 50 ns; sig_in <= "0011101111111101"; -- 0.468655
        wait for 50 ns; sig_in <= "0011001111001110"; -- 0.404711
        wait for 50 ns; sig_in <= "0010011111001001"; -- 0.310835
        wait for 50 ns; sig_in <= "0001100011001101"; -- 0.193766
        wait for 50 ns; sig_in <= "0000011111110001"; -- 0.062040
        wait for 50 ns; sig_in <= "1111011001110011"; -- -0.074610
        wait for 50 ns; sig_in <= "1110010110100011"; -- -0.205974
        wait for 50 ns; sig_in <= "1101011011000101"; -- -0.322120
        wait for 50 ns; sig_in <= "1100101011111101"; -- -0.414159
        wait for 50 ns; sig_in <= "1100001100110101"; -- -0.474932
        wait for 50 ns; sig_in <= "1100000000001110"; -- -0.499587
        wait for 50 ns; sig_in <= "1100000111001011"; -- -0.485989
        wait for 50 ns; sig_in <= "1100100001010100"; -- -0.434930
        wait for 50 ns; sig_in <= "1101001100110000"; -- -0.350109
        wait for 50 ns; sig_in <= "1110000110001101"; -- -0.237892
        wait for 50 ns; sig_in <= "1111001001010010"; -- -0.106859
        wait for 50 ns; sig_in <= "0000010000110100"; -- 0.032840
        wait for 50 ns; sig_in <= "0001010111001011"; -- 0.170257
        wait for 50 ns; sig_in <= "0010010110110010"; -- 0.294503
        wait for 50 ns; sig_in <= "0011001010100100"; -- 0.395617
        wait for 50 ns; sig_in <= "0011101110010001"; -- 0.465373
        wait for 50 ns; sig_in <= "0011111110111110"; -- 0.497972
        wait for 50 ns; sig_in <= "0011111011001010"; -- 0.490544
        wait for 50 ns; sig_in <= "0011100011000010"; -- 0.443428
        wait for 50 ns; sig_in <= "0010111000011011"; -- 0.360190
        wait for 50 ns; sig_in <= "0001111110101010"; -- 0.247389
        wait for 50 ns; sig_in <= "0000111010011010"; -- 0.114075
        wait for 50 ns; sig_in <= "1111110001001101"; -- -0.028911
        wait for 50 ns; sig_in <= "1110101001000100"; -- -0.169812
        wait for 50 ns; sig_in <= "1101100111111111"; -- -0.296913
        wait for 50 ns; sig_in <= "1100110011011100"; -- -0.399529
        wait for 50 ns; sig_in <= "1100001111111011"; -- -0.468907
        wait for 50 ns; sig_in <= "1100000000100001"; -- -0.498997
        wait for 50 ns; sig_in <= "1100000110101010"; -- -0.487007
        wait for 50 ns; sig_in <= "1100100001111101"; -- -0.433684
        wait for 50 ns; sig_in <= "1101010000001111"; -- -0.343307
        wait for 50 ns; sig_in <= "1110001101101001"; -- -0.223372
        wait for 50 ns; sig_in <= "1111010101000000"; -- -0.083998
        wait for 50 ns; sig_in <= "0000100000001110"; -- 0.062913
        wait for 50 ns; sig_in <= "0001101000110011"; -- 0.204678
        wait for 50 ns; sig_in <= "0010101000011010"; -- 0.328926
        wait for 50 ns; sig_in <= "0011011001011100"; -- 0.424690
        wait for 50 ns; sig_in <= "0011110111100000"; -- 0.483386
        wait for 50 ns; sig_in <= "0011111111110011"; -- 0.499608
        wait for 50 ns; sig_in <= "0011110001011111"; -- 0.471656
        wait for 50 ns; sig_in <= "0011001101101100"; -- 0.401736
        wait for 50 ns; sig_in <= "0010010111011110"; -- 0.295828
        wait for 50 ns; sig_in <= "0001010011100100"; -- 0.163198
        wait for 50 ns; sig_in <= "0000001000000000"; -- 0.015616
        wait for 50 ns; sig_in <= "1110111011100100"; -- -0.133677
        wait for 50 ns; sig_in <= "1101110101001011"; -- -0.271144
        wait for 50 ns; sig_in <= "1100111011010011"; -- -0.384188
        wait for 50 ns; sig_in <= "1100010011010011"; -- -0.462316
        wait for 50 ns; sig_in <= "1100000000111101"; -- -0.498138
        wait for 50 ns; sig_in <= "1100000110000110"; -- -0.488090
        wait for 50 ns; sig_in <= "1100100010011001"; -- -0.432821
        wait for 50 ns; sig_in <= "1101010011010111"; -- -0.337197
        wait for 50 ns; sig_in <= "1110010100100010"; -- -0.209900
        wait for 50 ns; sig_in <= "1111011111111010"; -- -0.062673
        wait for 50 ns; sig_in <= "0000101110011110"; -- 0.090745
        wait for 50 ns; sig_in <= "0001111000110010"; -- 0.235890
        wait for 50 ns; sig_in <= "0010110111110010"; -- 0.358938
        wait for 50 ns; sig_in <= "0011100101011001"; -- 0.448030
        wait for 50 ns; sig_in <= "0011111101001010"; -- 0.494439
        wait for 50 ns; sig_in <= "0011111100101001"; -- 0.493450
        wait for 50 ns; sig_in <= "0011100011110010"; -- 0.444876
        wait for 50 ns; sig_in <= "0010110100110100"; -- 0.353136
        wait for 50 ns; sig_in <= "0001110100001011"; -- 0.226890
        wait for 50 ns; sig_in <= "0000101000000100"; -- 0.078256
        wait for 50 ns; sig_in <= "1111010111111001"; -- -0.078334
        wait for 50 ns; sig_in <= "1110001011100001"; -- -0.227521
        wait for 50 ns; sig_in <= "1101001010011111"; -- -0.354526
        wait for 50 ns; sig_in <= "1100011011010101"; -- -0.446623
        wait for 50 ns; sig_in <= "1100000010110110"; -- -0.494438
        wait for 50 ns; sig_in <= "1100000011101000"; -- -0.492933
        wait for 50 ns; sig_in <= "1100011101101110"; -- -0.441968
        wait for 50 ns; sig_in <= "1101001110101010"; -- -0.346389
        wait for 50 ns; sig_in <= "1110010001100111"; -- -0.215600
        wait for 50 ns; sig_in <= "1111011111111010"; -- -0.062676
        wait for 50 ns; sig_in <= "0000110001101000"; -- 0.096926
        wait for 50 ns; sig_in <= "0001111110011011"; -- 0.246914
        wait for 50 ns; sig_in <= "0010111110011000"; -- 0.371825
        wait for 50 ns; sig_in <= "0011101010110101"; -- 0.458635
        wait for 50 ns; sig_in <= "0011111111000011"; -- 0.498138
        wait for 50 ns; sig_in <= "0011111000110100"; -- 0.485955
        wait for 50 ns; sig_in <= "0011011000100111"; -- 0.423061
        wait for 50 ns; sig_in <= "0010100001101011"; -- 0.315752
        wait for 50 ns; sig_in <= "0001011001101000"; -- 0.175053
        wait for 50 ns; sig_in <= "0000001000000000"; -- 0.015622
        wait for 50 ns; sig_in <= "1110110101011000"; -- -0.145760
        wait for 50 ns; sig_in <= "1101101010100010"; -- -0.291945
        wait for 50 ns; sig_in <= "1100101111100000"; -- -0.407241
        wait for 50 ns; sig_in <= "1100001010101100"; -- -0.479121
        wait for 50 ns; sig_in <= "1100000000001101"; -- -0.499608
        wait for 50 ns; sig_in <= "1100010001010100"; -- -0.466202
        wait for 50 ns; sig_in <= "1100111100010100"; -- -0.382217
        wait for 50 ns; sig_in <= "1101111100101011"; -- -0.256507
        wait for 50 ns; sig_in <= "1111001011011111"; -- -0.102562
        wait for 50 ns; sig_in <= "0000100000001101"; -- 0.062904
        wait for 50 ns; sig_in <= "0001110001100010"; -- 0.221751
        wait for 50 ns; sig_in <= "0010110110011111"; -- 0.356404
        wait for 50 ns; sig_in <= "0011100111010101"; -- 0.451803
        wait for 50 ns; sig_in <= "0011111110100010"; -- 0.497117
        wait for 50 ns; sig_in <= "0011111001010110"; -- 0.487010
        wait for 50 ns; sig_in <= "0011011000001110"; -- 0.422306
        wait for 50 ns; sig_in <= "0010011110101110"; -- 0.309984
        wait for 50 ns; sig_in <= "0001010011001100"; -- 0.162463
        wait for 50 ns; sig_in <= "1111111110000110"; -- -0.003732
        wait for 50 ns; sig_in <= "1110101001000100"; -- -0.169800
        wait for 50 ns; sig_in <= "1101011101110100"; -- -0.316781
        wait for 50 ns; sig_in <= "1100100101000000"; -- -0.427729
        wait for 50 ns; sig_in <= "1100000101010010"; -- -0.489688
        wait for 50 ns; sig_in <= "1100000010011100"; -- -0.495240
        wait for 50 ns; sig_in <= "1100011100111110"; -- -0.443434
        wait for 50 ns; sig_in <= "1101010001111011"; -- -0.339983
        wait for 50 ns; sig_in <= "1110011011010011"; -- -0.196680
        wait for 50 ns; sig_in <= "1111110000100110"; -- -0.030091
        wait for 50 ns; sig_in <= "0001000111110110"; -- 0.140327
        wait for 50 ns; sig_in <= "0010010110110010"; -- 0.294491
        wait for 50 ns; sig_in <= "0011010100000000"; -- 0.414061
        wait for 50 ns; sig_in <= "0011111000001001"; -- 0.484646
        wait for 50 ns; sig_in <= "0011111110110000"; -- 0.497564
        wait for 50 ns; sig_in <= "0011100110111001"; -- 0.450963
        wait for 50 ns; sig_in <= "0010110011010001"; -- 0.350121
        wait for 50 ns; sig_in <= "0001101001111100"; -- 0.206905
        wait for 50 ns; sig_in <= "0000010011101011"; -- 0.038415
        wait for 50 ns; sig_in <= "1110111010110111"; -- -0.135029
        wait for 50 ns; sig_in <= "1101101010010101"; -- -0.292323
        wait for 50 ns; sig_in <= "1100101011111101"; -- -0.414149
        wait for 50 ns; sig_in <= "1100000111011111"; -- -0.485372
        wait for 50 ns; sig_in <= "1100000001100100"; -- -0.496957
        wait for 50 ns; sig_in <= "1100011011000100"; -- -0.447157
        wait for 50 ns; sig_in <= "1101010000111111"; -- -0.341828
        wait for 50 ns; sig_in <= "1110011100110010"; -- -0.193785
        wait for 50 ns; sig_in <= "1111110101000110"; -- -0.021292
        wait for 50 ns; sig_in <= "0001001110111100"; -- 0.154161
        wait for 50 ns; sig_in <= "0010011110111111"; -- 0.310526
        wait for 50 ns; sig_in <= "0011011011001000"; -- 0.427971
        wait for 50 ns; sig_in <= "0011111011100111"; -- 0.491421
        wait for 50 ns; sig_in <= "0011111100001011"; -- 0.492534
        wait for 50 ns; sig_in <= "0011011100100110"; -- 0.430845
        wait for 50 ns; sig_in <= "0010100000101111"; -- 0.313925
        wait for 50 ns; sig_in <= "0001010000001000"; -- 0.156502
        wait for 50 ns; sig_in <= "1111110101000100"; -- -0.021347
        wait for 50 ns; sig_in <= "1110011011010001"; -- -0.196733
        wait for 50 ns; sig_in <= "1101001110011001"; -- -0.346889
        wait for 50 ns; sig_in <= "1100011000100000"; -- -0.452136
        wait for 50 ns; sig_in <= "1100000000110001"; -- -0.498498
        wait for 50 ns; sig_in <= "1100001010011101"; -- -0.479596
        wait for 50 ns; sig_in <= "1100110100011100"; -- -0.397586
        wait for 50 ns; sig_in <= "1101111001010111"; -- -0.262970
        wait for 50 ns; sig_in <= "1111010000001110"; -- -0.093310
        wait for 50 ns; sig_in <= "0000101101100101"; -- 0.089027
        wait for 50 ns; sig_in <= "0010000101000001"; -- 0.259793
        wait for 50 ns; sig_in <= "0011001010110011"; -- 0.396084
        wait for 50 ns; sig_in <= "0011110101011110"; -- 0.479432
        wait for 50 ns; sig_in <= "0011111111001010"; -- 0.498344
        wait for 50 ns; sig_in <= "0011100110011000"; -- 0.449941
        wait for 50 ns; sig_in <= "0010101110010100"; -- 0.340450
        wait for 50 ns; sig_in <= "0001011110011101"; -- 0.184464
        wait for 50 ns; sig_in <= "0000000001100100"; -- 0.003046
        wait for 50 ns; sig_in <= "1110100100010100"; -- -0.179083
        wait for 50 ns; sig_in <= "1101010011100001"; -- -0.336896
        wait for 50 ns; sig_in <= "1100011010010111"; -- -0.448510
        wait for 50 ns; sig_in <= "1100000000111001"; -- -0.498257
        wait for 50 ns; sig_in <= "1100001010110011"; -- -0.478924
        wait for 50 ns; sig_in <= "1100110110110111"; -- -0.392864
        wait for 50 ns; sig_in <= "1101111111000110"; -- -0.251773
        wait for 50 ns; sig_in <= "1111011001100001"; -- -0.075163
        wait for 50 ns; sig_in <= "0000111001100000"; -- 0.112301
        wait for 50 ns; sig_in <= "0010010001100001"; -- 0.284215
        wait for 50 ns; sig_in <= "0011010101000101"; -- 0.416162
        wait for 50 ns; sig_in <= "0011111010011110"; -- 0.489203
        wait for 50 ns; sig_in <= "0011111100001111"; -- 0.492643
        wait for 50 ns; sig_in <= "0011011001111100"; -- 0.425650
        wait for 50 ns; sig_in <= "0010011000010100"; -- 0.297493
        wait for 50 ns; sig_in <= "0001000000101011"; -- 0.126321
        wait for 50 ns; sig_in <= "1111011111100100"; -- -0.063358
        wait for 50 ns; sig_in <= "1110000010111111"; -- -0.244157
        wait for 50 ns; sig_in <= "1100111000011101"; -- -0.389755
        wait for 50 ns; sig_in <= "1100001010111000"; -- -0.478755
        wait for 50 ns; sig_in <= "1100000001000110"; -- -0.497866
        wait for 50 ns; sig_in <= "1100011100101101"; -- -0.443948
        wait for 50 ns; sig_in <= "1101011001110100"; -- -0.324590
        wait for 50 ns; sig_in <= "1110101111100100"; -- -0.157108
        wait for 50 ns; sig_in <= "0000010001010111"; -- 0.033911
        wait for 50 ns; sig_in <= "0001110000101111"; -- 0.220184
        wait for 50 ns; sig_in <= "0010111111011100"; -- 0.373910
        wait for 50 ns; sig_in <= "0011110001101000"; -- 0.471937
        wait for 50 ns; sig_in <= "0011111111101001"; -- 0.499287
        wait for 50 ns; sig_in <= "0011100111001011"; -- 0.451511
        wait for 50 ns; sig_in <= "0010101011110001"; -- 0.335467
        wait for 50 ns; sig_in <= "0001010110001111"; -- 0.168419
        wait for 50 ns; sig_in <= "1111110011011110"; -- -0.024482
        wait for 50 ns; sig_in <= "1110010010011101"; -- -0.213944
        wait for 50 ns; sig_in <= "1101000010000100"; -- -0.370969
        wait for 50 ns; sig_in <= "1100001110101100"; -- -0.471309
        wait for 50 ns; sig_in <= "1100000000011000"; -- -0.499254
        wait for 50 ns; sig_in <= "1100011001100001"; -- -0.450150
        wait for 50 ns; sig_in <= "1101010110011010"; -- -0.331246
        wait for 50 ns; sig_in <= "1110101101101110"; -- -0.160692
        wait for 50 ns; sig_in <= "0000010010000000"; -- 0.035164
        wait for 50 ns; sig_in <= "0001110011101000"; -- 0.225816
        wait for 50 ns; sig_in <= "0011000011010000"; -- 0.381335
        wait for 50 ns; sig_in <= "0011110100010001"; -- 0.477089
        wait for 50 ns; sig_in <= "0011111110110100"; -- 0.497688
        wait for 50 ns; sig_in <= "0011100001000010"; -- 0.439527
        wait for 50 ns; sig_in <= "0010011111011111"; -- 0.311479
        wait for 50 ns; sig_in <= "0001000100011011"; -- 0.133622
        wait for 50 ns; sig_in <= "1111011110010010"; -- -0.065849
        wait for 50 ns; sig_in <= "1101111101011010"; -- -0.255061
        wait for 50 ns; sig_in <= "1100110001011001"; -- -0.403543
        wait for 50 ns; sig_in <= "1100000110100101"; -- -0.487162
        wait for 50 ns; sig_in <= "1100000100000011"; -- -0.492096
        wait for 50 ns; sig_in <= "1100101010011010"; -- -0.417186
        wait for 50 ns; sig_in <= "1101110011100101"; -- -0.274264
        wait for 50 ns; sig_in <= "1111010011110010"; -- -0.086355
        wait for 50 ns; sig_in <= "0000111011011000"; -- 0.115969
        wait for 50 ns; sig_in <= "0010011001010111"; -- 0.299540
        wait for 50 ns; sig_in <= "0011011110001110"; -- 0.434025
        wait for 50 ns; sig_in <= "0011111110011101"; -- 0.496978
        wait for 50 ns; sig_in <= "0011110100100011"; -- 0.477642
        wait for 50 ns; sig_in <= "0011000001111111"; -- 0.378863
        wait for 50 ns; sig_in <= "0001101110111111"; -- 0.216760
        wait for 50 ns; sig_in <= "0000001001010011"; -- 0.018164
        wait for 50 ns; sig_in <= "1110100001111010"; -- -0.183765
        wait for 50 ns; sig_in <= "1101001010001101"; -- -0.355060
        wait for 50 ns; sig_in <= "1100010001000100"; -- -0.466672
        wait for 50 ns; sig_in <= "1100000000010010"; -- -0.499439
        wait for 50 ns; sig_in <= "1100011010111010"; -- -0.447447
        wait for 50 ns; sig_in <= "1101011100100101"; -- -0.319177
        wait for 50 ns; sig_in <= "1110111010010001"; -- -0.136203
        wait for 50 ns; sig_in <= "0000100100000010"; -- 0.070366
        wait for 50 ns; sig_in <= "0010000111110000"; -- 0.265138
        wait for 50 ns; sig_in <= "0011010100001110"; -- 0.414490
        wait for 50 ns; sig_in <= "0011111100000111"; -- 0.492404
        wait for 50 ns; sig_in <= "0011111000010110"; -- 0.485059
        wait for 50 ns; sig_in <= "0011001001011010"; -- 0.393359
        wait for 50 ns; sig_in <= "0001110111010001"; -- 0.232928
        wait for 50 ns; sig_in <= "0000010000001001"; -- 0.031529
        wait for 50 ns; sig_in <= "1110100110000011"; -- -0.175684
        wait for 50 ns; sig_in <= "1101001011101001"; -- -0.352276
        wait for 50 ns; sig_in <= "1100010000111011"; -- -0.466952
        wait for 50 ns; sig_in <= "1100000000011100"; -- -0.499147
        wait for 50 ns; sig_in <= "1100011101010011"; -- -0.442790
        wait for 50 ns; sig_in <= "1101100010100011"; -- -0.307529
        wait for 50 ns; sig_in <= "1111000100000000"; -- -0.117176
        wait for 50 ns; sig_in <= "0000110000010110"; -- 0.094423
        wait for 50 ns; sig_in <= "0010010100001010"; -- 0.289359
        wait for 50 ns; sig_in <= "0011011101011011"; -- 0.432451
        wait for 50 ns; sig_in <= "0011111110110010"; -- 0.497629
        wait for 50 ns; sig_in <= "0011110010000011"; -- 0.472755
        wait for 50 ns; sig_in <= "0010111001010101"; -- 0.361961
        wait for 50 ns; sig_in <= "0001011110110000"; -- 0.185067
        wait for 50 ns; sig_in <= "1111110010110000"; -- -0.025885
        wait for 50 ns; sig_in <= "1110001001000001"; -- -0.232382
        wait for 50 ns; sig_in <= "1100110101000001"; -- -0.396456
        wait for 50 ns; sig_in <= "1100000110010011"; -- -0.487687
        wait for 50 ns; sig_in <= "1100000101101100"; -- -0.488903
        wait for 50 ns; sig_in <= "1100110011011101"; -- -0.399500
        wait for 50 ns; sig_in <= "1110000111010100"; -- -0.235713
        wait for 50 ns; sig_in <= "1111110001110010"; -- -0.027763
        wait for 50 ns; sig_in <= "0001011111000100"; -- 0.185659
        wait for 50 ns; sig_in <= "0010111010101010"; -- 0.364562
        wait for 50 ns; sig_in <= "0011110011010010"; -- 0.475163
        wait for 50 ns; sig_in <= "0011111110001000"; -- 0.496323
        wait for 50 ns; sig_in <= "0011011000111011"; -- 0.423666
        wait for 50 ns; sig_in <= "0010001010100010"; -- 0.270578
        wait for 50 ns; sig_in <= "0000100001101101"; -- 0.065834
        wait for 50 ns; sig_in <= "1110110010010100"; -- -0.151738
        wait for 50 ns; sig_in <= "1101010001101000"; -- -0.340584
        wait for 50 ns; sig_in <= "1100010010001111"; -- -0.464371
        wait for 50 ns; sig_in <= "1100000000100000"; -- -0.499024
        wait for 50 ns; sig_in <= "1100100000000000"; -- -0.437492
        wait for 50 ns; sig_in <= "1101101010110111"; -- -0.291276
        wait for 50 ns; sig_in <= "1111010010110000"; -- -0.088382
        wait for 50 ns; sig_in <= "0001000011100100"; -- 0.131967
        wait for 50 ns; sig_in <= "0010100111010111"; -- 0.326873
        wait for 50 ns; sig_in <= "0011101010100100"; -- 0.458117
        wait for 50 ns; sig_in <= "0011111111110110"; -- 0.499703
        wait for 50 ns; sig_in <= "0011100010110111"; -- 0.443085
        wait for 50 ns; sig_in <= "0010011001000111"; -- 0.299027
        wait for 50 ns; sig_in <= "0000110000111110"; -- 0.095655
        wait for 50 ns; sig_in <= "1110111111000000"; -- -0.126948
        wait for 50 ns; sig_in <= "1101011001110011"; -- -0.324603
        wait for 50 ns; sig_in <= "1100010101100111"; -- -0.457801
        wait for 50 ns; sig_in <= "1100000000001011"; -- -0.499652
        wait for 50 ns; sig_in <= "1100011110000000"; -- -0.441397
        wait for 50 ns; sig_in <= "1101101001010011"; -- -0.294340
        wait for 50 ns; sig_in <= "1111010011000100"; -- -0.087766
        wait for 50 ns; sig_in <= "0001000110000011"; -- 0.136815
        wait for 50 ns; sig_in <= "0010101010111111"; -- 0.333958
        wait for 50 ns; sig_in <= "0011101101010100"; -- 0.463489
        wait for 50 ns; sig_in <= "0011111111010111"; -- 0.498741
        wait for 50 ns; sig_in <= "0011011101010000"; -- 0.432133
        wait for 50 ns; sig_in <= "0010001101110010"; -- 0.276905
        wait for 50 ns; sig_in <= "0000100001000101"; -- 0.064591
        wait for 50 ns; sig_in <= "1110101101011011"; -- -0.161299
        wait for 50 ns; sig_in <= "1101001010101011"; -- -0.354161
        wait for 50 ns; sig_in <= "1100001101010111"; -- -0.473921
        wait for 50 ns; sig_in <= "1100000010010110"; -- -0.495417
        wait for 50 ns; sig_in <= "1100101100001001"; -- -0.413782
        wait for 50 ns; sig_in <= "1110000010001110"; -- -0.245654
        wait for 50 ns; sig_in <= "1111110010110000"; -- -0.025886
        wait for 50 ns; sig_in <= "0001100110001100"; -- 0.199593
        wait for 50 ns; sig_in <= "0011000100010010"; -- 0.383349
        wait for 50 ns; sig_in <= "0011111001000100"; -- 0.486439
        wait for 50 ns; sig_in <= "0011111001001101"; -- 0.486732
        wait for 50 ns; sig_in <= "0011000100011111"; -- 0.383762
        wait for 50 ns; sig_in <= "0001100101111010"; -- 0.199029
        wait for 50 ns; sig_in <= "1111110001011110"; -- -0.028387
        wait for 50 ns; sig_in <= "1101111111111111"; -- -0.250016
        wait for 50 ns; sig_in <= "1100101001110101"; -- -0.418313
        wait for 50 ns; sig_in <= "1100000001100110"; -- -0.496889
        wait for 50 ns; sig_in <= "1100010000001010"; -- -0.468455
        wait for 50 ns; sig_in <= "1101010010100100"; -- -0.338742
        wait for 50 ns; sig_in <= "1110111010101001"; -- -0.135464
        wait for 50 ns; sig_in <= "0000110001111011"; -- 0.097497
        wait for 50 ns; sig_in <= "0010011110011110"; -- 0.309508
        wait for 50 ns; sig_in <= "0011101000100011"; -- 0.454183
        wait for 50 ns; sig_in <= "0011111111110010"; -- 0.499579
        wait for 50 ns; sig_in <= "0011011110111001"; -- 0.435347
        wait for 50 ns; sig_in <= "0010001100111010"; -- 0.275204
        wait for 50 ns; sig_in <= "0000011011101110"; -- 0.054127
        wait for 50 ns; sig_in <= "1110100100010000"; -- -0.179198
        wait for 50 ns; sig_in <= "1101000001000000"; -- -0.373053
        wait for 50 ns; sig_in <= "1100001000000111"; -- -0.484167
        wait for 50 ns; sig_in <= "1100000110011011"; -- -0.487444
        wait for 50 ns; sig_in <= "1100111100100011"; -- -0.381740
        wait for 50 ns; sig_in <= "1110011110100011"; -- -0.190335
        wait for 50 ns; sig_in <= "0000010110100100"; -- 0.044079
        wait for 50 ns; sig_in <= "0010001001101010"; -- 0.268845
        wait for 50 ns; sig_in <= "0011011101110001"; -- 0.433150
        wait for 50 ns; sig_in <= "0011111111110001"; -- 0.499551
        wait for 50 ns; sig_in <= "0011100111101111"; -- 0.452600
        wait for 50 ns; sig_in <= "0010011010111010"; -- 0.302557
        wait for 50 ns; sig_in <= "0000101010101001"; -- 0.083279
        wait for 50 ns; sig_in <= "1110110000011111"; -- -0.155318
        wait for 50 ns; sig_in <= "1101001000011010"; -- -0.358571
        wait for 50 ns; sig_in <= "1100001010011101"; -- -0.479599
        wait for 50 ns; sig_in <= "1100000101000010"; -- -0.490187
        wait for 50 ns; sig_in <= "1100111001100111"; -- -0.387474
        wait for 50 ns; sig_in <= "1110011100001111"; -- -0.194840
        wait for 50 ns; sig_in <= "0000010110001011"; -- 0.043292
        wait for 50 ns; sig_in <= "0010001011000101"; -- 0.271624
        wait for 50 ns; sig_in <= "0011011111101001"; -- 0.436797
        wait for 50 ns; sig_in <= "0011111111111101"; -- 0.499906
        wait for 50 ns; sig_in <= "0011100100001111"; -- 0.445761
        wait for 50 ns; sig_in <= "0010010010110001"; -- 0.286666
        wait for 50 ns; sig_in <= "0000011110100110"; -- 0.059763
        wait for 50 ns; sig_in <= "1110100011000011"; -- -0.181541
        wait for 50 ns; sig_in <= "1100111101011001"; -- -0.380089
        wait for 50 ns; sig_in <= "1100000101111000"; -- -0.488535
        wait for 50 ns; sig_in <= "1100001001111000"; -- -0.480706
        wait for 50 ns; sig_in <= "1101001000101100"; -- -0.358045
        wait for 50 ns; sig_in <= "1110110011011101"; -- -0.149503
        wait for 50 ns; sig_in <= "0000110000101111"; -- 0.095171
        wait for 50 ns; sig_in <= "0010100010011011"; -- 0.317227
        wait for 50 ns; sig_in <= "0011101101000100"; -- 0.463009
        wait for 50 ns; sig_in <= "0011111110011101"; -- 0.496979
        wait for 50 ns; sig_in <= "0011010010001011"; -- 0.410493
        wait for 50 ns; sig_in <= "0001110010110000"; -- 0.224134
        wait for 50 ns; sig_in <= "1111110111010001"; -- -0.017054
        wait for 50 ns; sig_in <= "1101111101110001"; -- -0.254354
        wait for 50 ns; sig_in <= "1100100100000001"; -- -0.429646
        wait for 50 ns; sig_in <= "1100000000001011"; -- -0.499674
        wait for 50 ns; sig_in <= "1100011011001110"; -- -0.446827
        wait for 50 ns; sig_in <= "1101101110110000"; -- -0.283696
        wait for 50 ns; sig_in <= "1111100110010010"; -- -0.050225
        wait for 50 ns; sig_in <= "0001100100010101"; -- 0.195965
        wait for 50 ns; sig_in <= "0011001001100110"; -- 0.393738
        wait for 50 ns; sig_in <= "0011111100110000"; -- 0.493655
        wait for 50 ns; sig_in <= "0011110000110110"; -- 0.470411
        wait for 50 ns; sig_in <= "0010101000101001"; -- 0.329385
        wait for 50 ns; sig_in <= "0000110110000010"; -- 0.105543
        wait for 50 ns; sig_in <= "1110110101101101"; -- -0.145101
        wait for 50 ns; sig_in <= "1101000111111110"; -- -0.359441
        wait for 50 ns; sig_in <= "1100001000101000"; -- -0.483167
        wait for 50 ns; sig_in <= "1100000111111000"; -- -0.484605
        wait for 50 ns; sig_in <= "1101000110001011"; -- -0.362957
        wait for 50 ns; sig_in <= "1110110011110101"; -- -0.148758
        wait for 50 ns; sig_in <= "0000110101000100"; -- 0.103649
        wait for 50 ns; sig_in <= "0010101000111000"; -- 0.329821
        wait for 50 ns; sig_in <= "0011110001011111"; -- 0.471661
        wait for 50 ns; sig_in <= "0011111100000111"; -- 0.492407
        wait for 50 ns; sig_in <= "0011000101110010"; -- 0.386285
        wait for 50 ns; sig_in <= "0001011100010011"; -- 0.180261
        wait for 50 ns; sig_in <= "1111011010110011"; -- -0.072667
        wait for 50 ns; sig_in <= "1101100010110100"; -- -0.307016
        wait for 50 ns; sig_in <= "1100010011100101"; -- -0.461748
        wait for 50 ns; sig_in <= "1100000001111100"; -- -0.496230
        wait for 50 ns; sig_in <= "1100110010101011"; -- -0.401028
        wait for 50 ns; sig_in <= "1110011001010010"; -- -0.200634
        wait for 50 ns; sig_in <= "0000011010111110"; -- 0.052679
        wait for 50 ns; sig_in <= "0010010101101101"; -- 0.292403
        wait for 50 ns; sig_in <= "0011101001000101"; -- 0.455222
        wait for 50 ns; sig_in <= "0011111110111000"; -- 0.497797
        wait for 50 ns; sig_in <= "0011010001000111"; -- 0.408421
        wait for 50 ns; sig_in <= "0001101011101110"; -- 0.210393
        wait for 50 ns; sig_in <= "1111101001100001"; -- -0.043905
        wait for 50 ns; sig_in <= "1101101101001100"; -- -0.286756
        wait for 50 ns; sig_in <= "1100011000000000"; -- -0.453115
        wait for 50 ns; sig_in <= "1100000000111111"; -- -0.498082
        wait for 50 ns; sig_in <= "1100101110100001"; -- -0.409147
        wait for 50 ns; sig_in <= "1110010100100101"; -- -0.209823
        wait for 50 ns; sig_in <= "0000010111110001"; -- 0.046412
        wait for 50 ns; sig_in <= "0010010100101010"; -- 0.290354
        wait for 50 ns; sig_in <= "0011101001010110"; -- 0.455740
        wait for 50 ns; sig_in <= "0011111110101000"; -- 0.497300
        wait for 50 ns; sig_in <= "0011001110011111"; -- 0.403275
        wait for 50 ns; sig_in <= "0001100101110110"; -- 0.198907
        wait for 50 ns; sig_in <= "1111100001001100"; -- -0.060181
        wait for 50 ns; sig_in <= "1101100100110111"; -- -0.303021
        wait for 50 ns; sig_in <= "1100010011000110"; -- -0.462706
        wait for 50 ns; sig_in <= "1100000010100111"; -- -0.494896
        wait for 50 ns; sig_in <= "1100111000001100"; -- -0.390256
        wait for 50 ns; sig_in <= "1110100101001101"; -- -0.177329
        wait for 50 ns; sig_in <= "0000101011100100"; -- 0.085093
        wait for 50 ns; sig_in <= "0010100101111100"; -- 0.324099
        wait for 50 ns; sig_in <= "0011110010001000"; -- 0.472899
        wait for 50 ns; sig_in <= "0011111010101010"; -- 0.489561
        wait for 50 ns; sig_in <= "0010111100111010"; -- 0.368970
        wait for 50 ns; sig_in <= "0001001010000001"; -- 0.144555
        wait for 50 ns; sig_in <= "1111000010001001"; -- -0.120815
        wait for 50 ns; sig_in <= "1101001011100110"; -- -0.352357
        wait for 50 ns; sig_in <= "1100000111111110"; -- -0.484435
        wait for 50 ns; sig_in <= "1100001010101000"; -- -0.479256
        wait for 50 ns; sig_in <= "1101010011000010"; -- -0.337836
        wait for 50 ns; sig_in <= "1111001100110011"; -- -0.100012
        wait for 50 ns; sig_in <= "0001010101010100"; -- 0.166620
        wait for 50 ns; sig_in <= "0011000101100011"; -- 0.385844
        wait for 50 ns; sig_in <= "0011111101001111"; -- 0.494613
        wait for 50 ns; sig_in <= "0011101100001100"; -- 0.461289
        wait for 50 ns; sig_in <= "0010010111000011"; -- 0.295005
        wait for 50 ns; sig_in <= "0000010110001100"; -- 0.043347
        wait for 50 ns; sig_in <= "1110001110110010"; -- -0.221121
        wait for 50 ns; sig_in <= "1100101000000101"; -- -0.421712
        wait for 50 ns; sig_in <= "1100000000000100"; -- -0.499890
        wait for 50 ns; sig_in <= "1100100010100101"; -- -0.432468
        wait for 50 ns; sig_in <= "1110000101110100"; -- -0.238661
        wait for 50 ns; sig_in <= "0000001100111010"; -- 0.025210
        wait for 50 ns; sig_in <= "0010010000010111"; -- 0.281957
        wait for 50 ns; sig_in <= "0011101001100000"; -- 0.456060
        wait for 50 ns; sig_in <= "0011111101111011"; -- 0.495937
        wait for 50 ns; sig_in <= "0011000111010111"; -- 0.389374
        wait for 50 ns; sig_in <= "0001010101101111"; -- 0.167438
        wait for 50 ns; sig_in <= "1111001010100011"; -- -0.104402
        wait for 50 ns; sig_in <= "1101001111000111"; -- -0.345476
        wait for 50 ns; sig_in <= "1100001000010001"; -- -0.483843
        wait for 50 ns; sig_in <= "1100001011010110"; -- -0.477844
        wait for 50 ns; sig_in <= "1101010111101010"; -- -0.328808
        wait for 50 ns; sig_in <= "1111010110100010"; -- -0.080980
        wait for 50 ns; sig_in <= "0001100010000001"; -- 0.191446
        wait for 50 ns; sig_in <= "0011010000000111"; -- 0.406462
        wait for 50 ns; sig_in <= "0011111111011110"; -- 0.498951
        wait for 50 ns; sig_in <= "0011100001100011"; -- 0.440527
        wait for 50 ns; sig_in <= "0001111111001100"; -- 0.248425
        wait for 50 ns; sig_in <= "1111110110000101"; -- -0.019388
        wait for 50 ns; sig_in <= "1101101111110110"; -- -0.281563
        wait for 50 ns; sig_in <= "1100010101011111"; -- -0.458036
        wait for 50 ns; sig_in <= "1100000010110011"; -- -0.494533
        wait for 50 ns; sig_in <= "1100111101101111"; -- -0.379414
        wait for 50 ns; sig_in <= "1110110100011100"; -- -0.147577
        wait for 50 ns; sig_in <= "0001000010100010"; -- 0.129946
        wait for 50 ns; sig_in <= "0010111100001111"; -- 0.367636
        wait for 50 ns; sig_in <= "0011111011110101"; -- 0.491837
        wait for 50 ns; sig_in <= "0011101101011010"; -- 0.463685
        wait for 50 ns; sig_in <= "0010010101001110"; -- 0.291443
        wait for 50 ns; sig_in <= "0000001110011111"; -- 0.028286
        wait for 50 ns; sig_in <= "1110000011000110"; -- -0.243959
        wait for 50 ns; sig_in <= "1100011110101000"; -- -0.440184
        wait for 50 ns; sig_in <= "1100000000101100"; -- -0.498654
        wait for 50 ns; sig_in <= "1100110010111010"; -- -0.400570
        wait for 50 ns; sig_in <= "1110100101101111"; -- -0.176313
        wait for 50 ns; sig_in <= "0000110101001001"; -- 0.103778
        wait for 50 ns; sig_in <= "0010110011111001"; -- 0.351340
        wait for 50 ns; sig_in <= "0011111001110010"; -- 0.487847
        wait for 50 ns; sig_in <= "0011110000011100"; -- 0.469615
        wait for 50 ns; sig_in <= "0010011010100111"; -- 0.301960
        wait for 50 ns; sig_in <= "0000010011011001"; -- 0.037869
        wait for 50 ns; sig_in <= "1110000101110110"; -- -0.238580
        wait for 50 ns; sig_in <= "1100011111010010"; -- -0.438907
        wait for 50 ns; sig_in <= "1100000000101110"; -- -0.498595
        wait for 50 ns; sig_in <= "1100110100001110"; -- -0.398015
        wait for 50 ns; sig_in <= "1110101001011100"; -- -0.169079
        wait for 50 ns; sig_in <= "0000111010101110"; -- 0.114680
        wait for 50 ns; sig_in <= "0010111001001001"; -- 0.361601
        wait for 50 ns; sig_in <= "0011111011101001"; -- 0.491493
        wait for 50 ns; sig_in <= "0011101100011100"; -- 0.461780
        wait for 50 ns; sig_in <= "0010010000001101"; -- 0.281646
        wait for 50 ns; sig_in <= "0000000100110101"; -- 0.009419
        wait for 50 ns; sig_in <= "1101110111101111"; -- -0.266150
        wait for 50 ns; sig_in <= "1100010111001011"; -- -0.454754
        wait for 50 ns; sig_in <= "1100000010111111"; -- -0.494181
        wait for 50 ns; sig_in <= "1101000010000011"; -- -0.370995
        wait for 50 ns; sig_in <= "1110111111110101"; -- -0.125329
        wait for 50 ns; sig_in <= "0001010010111100"; -- 0.161994
        wait for 50 ns; sig_in <= "0011001010101110"; -- 0.395938
        wait for 50 ns; sig_in <= "0011111111010101"; -- 0.498692
        wait for 50 ns; sig_in <= "0011011111000100"; -- 0.435679
        wait for 50 ns; sig_in <= "0001110100011011"; -- 0.227397
        wait for 50 ns; sig_in <= "1111100010110011"; -- -0.057030
        wait for 50 ns; sig_in <= "1101011010110100"; -- -0.322640
        wait for 50 ns; sig_in <= "1100001010000110"; -- -0.480293
        wait for 50 ns; sig_in <= "1100001011111100"; -- -0.476676
        wait for 50 ns; sig_in <= "1101011111111111"; -- -0.312520
        wait for 50 ns; sig_in <= "1111101010000111"; -- -0.042740
        wait for 50 ns; sig_in <= "0001111011110010"; -- 0.241748
        wait for 50 ns; sig_in <= "0011100011101000"; -- 0.444579
        wait for 50 ns; sig_in <= "0011111110010010"; -- 0.496629
        wait for 50 ns; sig_in <= "0011000010011011"; -- 0.379731
        wait for 50 ns; sig_in <= "0001000100001110"; -- 0.133240
        wait for 50 ns; sig_in <= "1110101110100110"; -- -0.159009
        wait for 50 ns; sig_in <= "1100110100101100"; -- -0.397086
        wait for 50 ns; sig_in <= "1100000000011100"; -- -0.499144
        wait for 50 ns; sig_in <= "1100100100000000"; -- -0.429688
        wait for 50 ns; sig_in <= "1110010011011001"; -- -0.212134
        wait for 50 ns; sig_in <= "0000101000011000"; -- 0.078854
        wait for 50 ns; sig_in <= "0010101111100010"; -- 0.342835
        wait for 50 ns; sig_in <= "0011111001111110"; -- 0.488221
        wait for 50 ns; sig_in <= "0011101101101010"; -- 0.464161
        wait for 50 ns; sig_in <= "0010001110100111"; -- 0.278525
        wait for 50 ns; sig_in <= "1111111101101111"; -- -0.004421
        wait for 50 ns; sig_in <= "1101101101100010"; -- -0.286083
        wait for 50 ns; sig_in <= "1100010000011110"; -- -0.467821
        wait for 50 ns; sig_in <= "1100000111011001"; -- -0.485569
        wait for 50 ns; sig_in <= "1101010101101101"; -- -0.332602
        wait for 50 ns; sig_in <= "1111100000000110"; -- -0.062311
        wait for 50 ns; sig_in <= "0001110101111000"; -- 0.230226
        wait for 50 ns; sig_in <= "0011100010000110"; -- 0.441586
        wait for 50 ns; sig_in <= "0011111110010001"; -- 0.496611
        wait for 50 ns; sig_in <= "0011000000001010"; -- 0.375298
        wait for 50 ns; sig_in <= "0000111101100110"; -- 0.120305
        wait for 50 ns; sig_in <= "1110100100111101"; -- -0.177822
        wait for 50 ns; sig_in <= "1100101100101101"; -- -0.412677
        wait for 50 ns; sig_in <= "1100000000000001"; -- -0.499984
        wait for 50 ns; sig_in <= "1100101111000111"; -- -0.407989
        wait for 50 ns; sig_in <= "1110101001010110"; -- -0.169241
        wait for 50 ns; sig_in <= "0001000010111010"; -- 0.130685
        wait for 50 ns; sig_in <= "0011000100011110"; -- 0.383713
        wait for 50 ns; sig_in <= "0011111111000101"; -- 0.498196
        wait for 50 ns; sig_in <= "0011011101010100"; -- 0.432246
        wait for 50 ns; sig_in <= "0001101011001010"; -- 0.209287
        wait for 50 ns; sig_in <= "1111010001111010"; -- -0.090016
        wait for 50 ns; sig_in <= "1101001001010101"; -- -0.356771
        wait for 50 ns; sig_in <= "1100000011010111"; -- -0.493445
        wait for 50 ns; sig_in <= "1100011001110010"; -- -0.449639
        wait for 50 ns; sig_in <= "1110000100101010"; -- -0.240899
        wait for 50 ns; sig_in <= "0000011100111101"; -- 0.056547
        wait for 50 ns; sig_in <= "0010101010101110"; -- 0.333437
        wait for 50 ns; sig_in <= "0011111001101001"; -- 0.487565
        wait for 50 ns; sig_in <= "0011101100010110"; -- 0.461606
        wait for 50 ns; sig_in <= "0010000111100000"; -- 0.264659
        wait for 50 ns; sig_in <= "1111110000010011"; -- -0.030677
        wait for 50 ns; sig_in <= "1101011110110010"; -- -0.314867
        wait for 50 ns; sig_in <= "1100001001001110"; -- -0.482000
        wait for 50 ns; sig_in <= "1100001111101100"; -- -0.469353
        wait for 50 ns; sig_in <= "1101110000000100"; -- -0.281143
        wait for 50 ns; sig_in <= "0000000110011101"; -- 0.012593
        wait for 50 ns; sig_in <= "0010011010100011"; -- 0.301859
        wait for 50 ns; sig_in <= "0011110100101001"; -- 0.477809
        wait for 50 ns; sig_in <= "0011110010100101"; -- 0.473796
        wait for 50 ns; sig_in <= "0010010100111010"; -- 0.290827
        wait for 50 ns; sig_in <= "1111111110110011"; -- -0.002362
        wait for 50 ns; sig_in <= "1101101001000000"; -- -0.294911
        wait for 50 ns; sig_in <= "1100001100011101"; -- -0.475674
        wait for 50 ns; sig_in <= "1100001100100010"; -- -0.475528
        wait for 50 ns; sig_in <= "1101101001011110"; -- -0.294020
        wait for 50 ns; sig_in <= "0000000000000000"; -- -0.000000
    end process;

END;
