package RTL_SVPackage;
   localparam CONST = 0;
endpackage // RTL_SVPackage
   
