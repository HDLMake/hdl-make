//                              -*- Mode: Verilog -*-
// Filename        : includeModuleSV.sv
// Description     : Included submodule
// Author          : Adrian Fiergolski
// Created On      : Thu Sep 18 10:51:41 2014
// Last Modified By: Adrian Fiergolski
// Last Modified On: Thu Sep 18 10:51:41 2014
// Update Count    : 0
// Status          : Unknown, Use with caution!

module includeModuleSV;


endmodule // includeModuleSV
